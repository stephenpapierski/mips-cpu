LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY dec5to32_tb IS
END dec5to32_tb;

ARCHITECTURE test OF dec5to32_tb IS
    SIGNAL i0 : STD_LOGIC_VECTOR(4 downto 0);
    SIGNAL w, q0, q1, q2, q3, q4, q5, q6, q7, q8, q9, q10, q11, q12, q13, q14, q15, q16, q17, q18, q19, q20, q21, q22, q23, q24, q25, q26, q27, q28, q29, q30, q31: STD_LOGIC;
BEGIN
    dec_0: ENTITY work.dec5to32(struct) PORT MAP (i0, w, q0, q1, q2, q3, q4, q5, q6, q7, q8, q9, q10, q11, q12, q13, q14, q15, q16, q17, q18, q19, q20, q21, q22, q23, q24, q25, q26, q27, q28, q29, q30, q31);

    PROCESS
	TYPE pattern_type IS RECORD
	    i0 : STD_LOGIC_VECTOR(4 downto 0);
	    w, q0, q1, q2, q3, q4, q5, q6, q7, q8, q9, q10, q11, q12, q13, q14, q15, q16, q17, q18, q19, q20, q21, q22, q23, q24, q25, q26, q27, q28, q29, q30, q31: STD_LOGIC;
	END RECORD;
	TYPE pattern_array IS ARRAY (NATURAL RANGE <>) OF pattern_type;
	CONSTANT patterns: pattern_array :=
	    (
         ("00000", '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("00001", '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("00010", '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("00011", '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("00100", '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("00101", '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("00110", '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("00111", '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("01000", '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("01001", '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("01010", '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("01011", '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("01100", '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("01101", '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("01110", '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("01111", '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("10000", '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("10001", '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("10010", '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("10011", '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("10100", '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("10101", '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("10110", '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("10111", '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("11000", '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("11001", '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("11010", '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("11011", '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("11100", '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("11101", '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("11110", '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("11111", '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         

         ("00000", '1', '1','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("00001", '1', '0','1', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("00010", '1', '0','0', '1', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("00011", '1', '0','0', '0', '1','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("00100", '1', '0','0', '0', '0','1', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("00101", '1', '0','0', '0', '0','0', '1', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("00110", '1', '0','0', '0', '0','0', '0', '1','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("00111", '1', '0','0', '0', '0','0', '0', '0','1', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("01000", '1', '0','0', '0', '0','0', '0', '0','0', '1', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("01001", '1', '0','0', '0', '0','0', '0', '0','0', '0', '1', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("01010", '1', '0','0', '0', '0','0', '0', '0','0', '0', '0', '1','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("01011", '1', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','1', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("01100", '1', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '1', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("01101", '1', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '1','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("01110", '1', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','1', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("01111", '1', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '1', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("10000", '1', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '1','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("10001", '1', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','1', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("10010", '1', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '1', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("10011", '1', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '1', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("10100", '1', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '1','0', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("10101", '1', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','1', '0', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("10110", '1', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '1', '0','0', '0', '0','0', '0', '0', '0', '0'),
         ("10111", '1', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '1','0', '0', '0','0', '0', '0', '0', '0'),
         ("11000", '1', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','1', '0', '0','0', '0', '0', '0', '0'),
         ("11001", '1', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '1', '0','0', '0', '0', '0', '0'),
         ("11010", '1', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '1','0', '0', '0', '0', '0'),
         ("11011", '1', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','1', '0', '0', '0', '0'),
         ("11100", '1', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '1', '0', '0', '0'),
         ("11101", '1', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '1', '0', '0'),
         ("11110", '1', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '1', '0'),
         ("11111", '1', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0','0', '0', '0','0', '0', '0','0', '0', '0', '0', '1')
     );
    BEGIN
      --  Check each pattern.
      for i in patterns'range loop
	  --  Set the inputs.
	  i0 <= patterns(i).i0;
	  w <= patterns(i).w;
	  q0 <= patterns(i).q0;
	  q1 <= patterns(i).q1;
	  q2 <= patterns(i).q2;
	  q3 <= patterns(i).q3;
	  q4 <= patterns(i).q4;
	  q5 <= patterns(i).q5;
	  q6 <= patterns(i).q6;
	  q7 <= patterns(i).q7;
	  q8 <= patterns(i).q8;
	  q9 <= patterns(i).q9;
	  q10 <= patterns(i).q10;
	  q11 <= patterns(i).q11;
	  q12 <= patterns(i).q12;
	  q13 <= patterns(i).q13;
	  q14 <= patterns(i).q14;
	  q15 <= patterns(i).q15;
	  q16 <= patterns(i).q16;
	  q17 <= patterns(i).q17;
	  q18 <= patterns(i).q18;
	  q19 <= patterns(i).q19;
	  q20 <= patterns(i).q20;
	  q21 <= patterns(i).q21;
	  q22 <= patterns(i).q22;
	  q23 <= patterns(i).q23;
	  q24 <= patterns(i).q24;
	  q25 <= patterns(i).q25;
	  q26 <= patterns(i).q26;
	  q27 <= patterns(i).q27;
	  q28 <= patterns(i).q28;
	  q29 <= patterns(i).q29;
	  q30 <= patterns(i).q30;
	  q31 <= patterns(i).q31;
	  --  Wait for the results.
	  wait for 1 ns;
	  --  Check the outputs.
	  --assert o1 = patterns(i).o
	  --  report "bad Behavior output value" severity error;
      end loop;
      assert false report "end of test" severity note;
      --  Wait forever; this will finish the simulation.
      wait;
    END PROCESS;
END test;
